/home/atreya/SSV/Tempus/tempus_labs/libs/MACRO/LEF/rom_512x16A.lef