../../../../libs/lef/FreePDK45_lib_v1.0.lef