../../../../libs/MACRO/LEF/ram_256X16A.lef