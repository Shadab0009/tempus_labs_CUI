../../../../libs/MACRO/LEF/pllclk.lef