../../../../libs/MACRO/LEF/rom_512x16A.lef