* Comment

.subckt ant in
.ends
