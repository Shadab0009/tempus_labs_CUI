module pllclk(refclk, vcop, vcom, clk1x, clk2x);
    input  refclk;
    output vcop;
    output vcom;
    output clk1x;
    output clk2x;
endmodule

