/home/atreya/SSV/Tempus/tempus_labs/libs/MACRO/LEF/pllclk.lef