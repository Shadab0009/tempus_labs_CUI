/home/atreya/SSV/Tempus/tempus_labs/libs/MACRO/LEF/ram_256X16A.lef